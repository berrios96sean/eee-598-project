module top (

    input clk,
    input rst,
    input x,
    output y
);



endmodule 
